library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
        tmp(0)  := "0100" & "0" & "00000100";   -- Desta posicao para baixo, é necessário acertar os valores
        tmp(1)  := "0101" & "1" & "00000001";
        tmp(2)  := "0100" & "0" & "00000011";
		  tmp(3)  := "0101" & "1" & "00000000";
        tmp(4)  := "0010" & "1" & "00000000";
		  tmp(5)  := "0010" & "1" & "00000000";
		  tmp(6)  := "0011" & "1" & "00000001";
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;